//ddfsdfsdf
//sdfsdfsdf



module 