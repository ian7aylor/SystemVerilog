//ddfsdfsdf
//sdfsdfsdf

